entity and2 is
port(
 in_port1 : in std_logic;
 in_port2 : in std_logic;

 out_port1 : out std_logic);
end and2;